module top #(
	parameter WIDTH = 16
)(
  // interface signals
  input  logic             clk,      // clock 
  input  logic             rst,      // reset
  output  logic            a0        // output signal
);

  // add stuff

endmodule